--------------------------------------------------------------------------------
--
--    Filename    : dmem_init.vhd
--    Entity      : dmem4
--    Input from  : dmem.bin
--    Description : Single Port Asynchronous Random Access (initialized) Data
--                  Memory with 4 write enable ports.
--    Author      : Tamar/Rene/Huib
--    Company     : Delft University of Technology
--
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.numeric_std.all;


ENTITY dmem4 IS
    GENERIC (
        WIDTH_g : POSITIVE := 32;
        ABITS_g : POSITIVE := 14
        );
    PORT (
        clk_i :  IN STD_LOGIC;
        ce_i  :  IN STD_LOGIC;
        adr_i :  IN STD_LOGIC_VECTOR (ABITS_g -1 DOWNTO 0);
        wre_i :  IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        dat_i :  IN STD_LOGIC_VECTOR (WIDTH_g -1 DOWNTO 0);
        dat_o : OUT STD_LOGIC_VECTOR (WIDTH_g -1 DOWNTO 0)
    );
END dmem4;


ARCHITECTURE arch OF dmem4 IS

    SIGNAL word_adr_s         : STD_LOGIC_VECTOR (  ABITS_g -3 DOWNTO 0);
    SIGNAL di0, di1, di2, di3 : STD_LOGIC_VECTOR (WIDTH_g/4 -1 DOWNTO 0);
    SIGNAL do0, do1, do2, do3 : STD_LOGIC_VECTOR (WIDTH_g/4 -1 DOWNTO 0);

    TYPE ram_type IS ARRAY (0 TO 2**(ABITS_g-2) -1) OF STD_LOGIC_VECTOR (WIDTH_g/4 -1 DOWNTO 0);

    SIGNAL ram0 : ram_type := (
         X"FF", X"00", X"FF", X"00", X"00", X"43", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00" );

    SIGNAL ram1 : ram_type := (
         X"FF", X"00", X"FF", X"00", X"00", X"00", X"00", X"00",
         X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00" );

    SIGNAL ram2 : ram_type := (
         X"FF", X"00", X"FF", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00" );

    SIGNAL ram3 : ram_type := (
         X"FF", X"00", X"FF", X"00", X"2C", X"00", X"00", X"00",
         X"0C", X"00", X"2C", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"14", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
         X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00" );


BEGIN


    word_adr_s <= adr_i(ABITS_g -1 DOWNTO 2);  -- convert to word-address

    do3   <= ram3(TO_INTEGER(UNSIGNED(word_adr_s)));
    do2   <= ram2(TO_INTEGER(UNSIGNED(word_adr_s)));
    do1   <= ram1(TO_INTEGER(UNSIGNED(word_adr_s)));
    do0   <= ram0(TO_INTEGER(UNSIGNED(word_adr_s)));
    dat_o <= do0 & do1 & do2 & do3;

    di3   <= dat_i(  WIDTH_g/4 -1 DOWNTO         0);
    di2   <= dat_i(  WIDTH_g/2 -1 DOWNTO   WIDTH_g/4);
    di1   <= dat_i(3*WIDTH_g/4 -1 DOWNTO   WIDTH_g/2);
    di0   <= dat_i(  WIDTH_g   -1 DOWNTO 3*WIDTH_g/4);

	PROCESS (clk_i)
	BEGIN
		IF FALLING_EDGE (clk_i) THEN
			IF (ce_i = '1') THEN
				IF (wre_i(0) = '1') THEN
	    			ram3(TO_INTEGER(UNSIGNED(word_adr_s))) <= di3;
	    		END IF;
				IF (wre_i(1) = '1') THEN
	    			ram2(TO_INTEGER(UNSIGNED(word_adr_s))) <= di2;
	    		END IF;
				IF (wre_i(2) = '1') THEN
	    			ram1(TO_INTEGER(UNSIGNED(word_adr_s))) <= di1;
	    		END IF;
				IF (wre_i(3) = '1') THEN
	    			ram0(TO_INTEGER(UNSIGNED(word_adr_s))) <= di0;
	    		END IF;
    		END IF;
   		END IF;
   	END PROCESS;

END ARCHITECTURE arch;

-- [EOF]
